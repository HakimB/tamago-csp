module tamago.example;

service Sudoku { 
 method void initGrille(int[] grille) {
id initGrille;
pre  (grille.length == 81) && 
(grille[0] != grille[1]) &&
(grille[0] != grille[2]) &&
(grille[0] != grille[3]) &&
(grille[0] != grille[4]) &&
(grille[0] != grille[5]) &&
(grille[0] != grille[6]) &&
(grille[0] != grille[7]) &&
(grille[0] != grille[8]) &&
(grille[1] != grille[2]) &&
(grille[1] != grille[3]) &&
(grille[1] != grille[4]) &&
(grille[1] != grille[5]) &&
(grille[1] != grille[6]) &&
(grille[1] != grille[7]) &&
(grille[1] != grille[8]) &&
(grille[2] != grille[3]) &&
(grille[2] != grille[4]) &&
(grille[2] != grille[5]) &&
(grille[2] != grille[6]) &&
(grille[2] != grille[7]) &&
(grille[2] != grille[8]) &&
(grille[3] != grille[4]) &&
(grille[3] != grille[5]) &&
(grille[3] != grille[6]) &&
(grille[3] != grille[7]) &&
(grille[3] != grille[8]) &&
(grille[4] != grille[5]) &&
(grille[4] != grille[6]) &&
(grille[4] != grille[7]) &&
(grille[4] != grille[8]) &&
(grille[5] != grille[6]) &&
(grille[5] != grille[7]) &&
(grille[5] != grille[8]) &&
(grille[6] != grille[7]) &&
(grille[6] != grille[8]) &&
(grille[7] != grille[8]) &&
(grille[9] != grille[10]) &&
(grille[9] != grille[11]) &&
(grille[9] != grille[12]) &&
(grille[9] != grille[13]) &&
(grille[9] != grille[14]) &&
(grille[9] != grille[15]) &&
(grille[9] != grille[16]) &&
(grille[9] != grille[17]) &&
(grille[10] != grille[11]) &&
(grille[10] != grille[12]) &&
(grille[10] != grille[13]) &&
(grille[10] != grille[14]) &&
(grille[10] != grille[15]) &&
(grille[10] != grille[16]) &&
(grille[10] != grille[17]) &&
(grille[11] != grille[12]) &&
(grille[11] != grille[13]) &&
(grille[11] != grille[14]) &&
(grille[11] != grille[15]) &&
(grille[11] != grille[16]) &&
(grille[11] != grille[17]) &&
(grille[12] != grille[13]) &&
(grille[12] != grille[14]) &&
(grille[12] != grille[15]) &&
(grille[12] != grille[16]) &&
(grille[12] != grille[17]) &&
(grille[13] != grille[14]) &&
(grille[13] != grille[15]) &&
(grille[13] != grille[16]) &&
(grille[13] != grille[17]) &&
(grille[14] != grille[15]) &&
(grille[14] != grille[16]) &&
(grille[14] != grille[17]) &&
(grille[15] != grille[16]) &&
(grille[15] != grille[17]) &&
(grille[16] != grille[17]) &&
(grille[18] != grille[19]) &&
(grille[18] != grille[20]) &&
(grille[18] != grille[21]) &&
(grille[18] != grille[22]) &&
(grille[18] != grille[23]) &&
(grille[18] != grille[24]) &&
(grille[18] != grille[25]) &&
(grille[18] != grille[26]) &&
(grille[19] != grille[20]) &&
(grille[19] != grille[21]) &&
(grille[19] != grille[22]) &&
(grille[19] != grille[23]) &&
(grille[19] != grille[24]) &&
(grille[19] != grille[25]) &&
(grille[19] != grille[26]) &&
(grille[20] != grille[21]) &&
(grille[20] != grille[22]) &&
(grille[20] != grille[23]) &&
(grille[20] != grille[24]) &&
(grille[20] != grille[25]) &&
(grille[20] != grille[26]) &&
(grille[21] != grille[22]) &&
(grille[21] != grille[23]) &&
(grille[21] != grille[24]) &&
(grille[21] != grille[25]) &&
(grille[21] != grille[26]) &&
(grille[22] != grille[23]) &&
(grille[22] != grille[24]) &&
(grille[22] != grille[25]) &&
(grille[22] != grille[26]) &&
(grille[23] != grille[24]) &&
(grille[23] != grille[25]) &&
(grille[23] != grille[26]) &&
(grille[24] != grille[25]) &&
(grille[24] != grille[26]) &&
(grille[25] != grille[26]) &&
(grille[27] != grille[28]) &&
(grille[27] != grille[29]) &&
(grille[27] != grille[30]) &&
(grille[27] != grille[31]) &&
(grille[27] != grille[32]) &&
(grille[27] != grille[33]) &&
(grille[27] != grille[34]) &&
(grille[27] != grille[35]) &&
(grille[28] != grille[29]) &&
(grille[28] != grille[30]) &&
(grille[28] != grille[31]) &&
(grille[28] != grille[32]) &&
(grille[28] != grille[33]) &&
(grille[28] != grille[34]) &&
(grille[28] != grille[35]) &&
(grille[29] != grille[30]) &&
(grille[29] != grille[31]) &&
(grille[29] != grille[32]) &&
(grille[29] != grille[33]) &&
(grille[29] != grille[34]) &&
(grille[29] != grille[35]) &&
(grille[30] != grille[31]) &&
(grille[30] != grille[32]) &&
(grille[30] != grille[33]) &&
(grille[30] != grille[34]) &&
(grille[30] != grille[35]) &&
(grille[31] != grille[32]) &&
(grille[31] != grille[33]) &&
(grille[31] != grille[34]) &&
(grille[31] != grille[35]) &&
(grille[32] != grille[33]) &&
(grille[32] != grille[34]) &&
(grille[32] != grille[35]) &&
(grille[33] != grille[34]) &&
(grille[33] != grille[35]) &&
(grille[34] != grille[35]) &&
(grille[36] != grille[37]) &&
(grille[36] != grille[38]) &&
(grille[36] != grille[39]) &&
(grille[36] != grille[40]) &&
(grille[36] != grille[41]) &&
(grille[36] != grille[42]) &&
(grille[36] != grille[43]) &&
(grille[36] != grille[44]) &&
(grille[37] != grille[38]) &&
(grille[37] != grille[39]) &&
(grille[37] != grille[40]) &&
(grille[37] != grille[41]) &&
(grille[37] != grille[42]) &&
(grille[37] != grille[43]) &&
(grille[37] != grille[44]) &&
(grille[38] != grille[39]) &&
(grille[38] != grille[40]) &&
(grille[38] != grille[41]) &&
(grille[38] != grille[42]) &&
(grille[38] != grille[43]) &&
(grille[38] != grille[44]) &&
(grille[39] != grille[40]) &&
(grille[39] != grille[41]) &&
(grille[39] != grille[42]) &&
(grille[39] != grille[43]) &&
(grille[39] != grille[44]) &&
(grille[40] != grille[41]) &&
(grille[40] != grille[42]) &&
(grille[40] != grille[43]) &&
(grille[40] != grille[44]) &&
(grille[41] != grille[42]) &&
(grille[41] != grille[43]) &&
(grille[41] != grille[44]) &&
(grille[42] != grille[43]) &&
(grille[42] != grille[44]) &&
(grille[43] != grille[44]) &&
(grille[45] != grille[46]) &&
(grille[45] != grille[47]) &&
(grille[45] != grille[48]) &&
(grille[45] != grille[49]) &&
(grille[45] != grille[50]) &&
(grille[45] != grille[51]) &&
(grille[45] != grille[52]) &&
(grille[45] != grille[53]) &&
(grille[46] != grille[47]) &&
(grille[46] != grille[48]) &&
(grille[46] != grille[49]) &&
(grille[46] != grille[50]) &&
(grille[46] != grille[51]) &&
(grille[46] != grille[52]) &&
(grille[46] != grille[53]) &&
(grille[47] != grille[48]) &&
(grille[47] != grille[49]) &&
(grille[47] != grille[50]) &&
(grille[47] != grille[51]) &&
(grille[47] != grille[52]) &&
(grille[47] != grille[53]) &&
(grille[48] != grille[49]) &&
(grille[48] != grille[50]) &&
(grille[48] != grille[51]) &&
(grille[48] != grille[52]) &&
(grille[48] != grille[53]) &&
(grille[49] != grille[50]) &&
(grille[49] != grille[51]) &&
(grille[49] != grille[52]) &&
(grille[49] != grille[53]) &&
(grille[50] != grille[51]) &&
(grille[50] != grille[52]) &&
(grille[50] != grille[53]) &&
(grille[51] != grille[52]) &&
(grille[51] != grille[53]) &&
(grille[52] != grille[53]) &&
(grille[54] != grille[55]) &&
(grille[54] != grille[56]) &&
(grille[54] != grille[57]) &&
(grille[54] != grille[58]) &&
(grille[54] != grille[59]) &&
(grille[54] != grille[60]) &&
(grille[54] != grille[61]) &&
(grille[54] != grille[62]) &&
(grille[55] != grille[56]) &&
(grille[55] != grille[57]) &&
(grille[55] != grille[58]) &&
(grille[55] != grille[59]) &&
(grille[55] != grille[60]) &&
(grille[55] != grille[61]) &&
(grille[55] != grille[62]) &&
(grille[56] != grille[57]) &&
(grille[56] != grille[58]) &&
(grille[56] != grille[59]) &&
(grille[56] != grille[60]) &&
(grille[56] != grille[61]) &&
(grille[56] != grille[62]) &&
(grille[57] != grille[58]) &&
(grille[57] != grille[59]) &&
(grille[57] != grille[60]) &&
(grille[57] != grille[61]) &&
(grille[57] != grille[62]) &&
(grille[58] != grille[59]) &&
(grille[58] != grille[60]) &&
(grille[58] != grille[61]) &&
(grille[58] != grille[62]) &&
(grille[59] != grille[60]) &&
(grille[59] != grille[61]) &&
(grille[59] != grille[62]) &&
(grille[60] != grille[61]) &&
(grille[60] != grille[62]) &&
(grille[61] != grille[62]) &&
(grille[63] != grille[64]) &&
(grille[63] != grille[65]) &&
(grille[63] != grille[66]) &&
(grille[63] != grille[67]) &&
(grille[63] != grille[68]) &&
(grille[63] != grille[69]) &&
(grille[63] != grille[70]) &&
(grille[63] != grille[71]) &&
(grille[64] != grille[65]) &&
(grille[64] != grille[66]) &&
(grille[64] != grille[67]) &&
(grille[64] != grille[68]) &&
(grille[64] != grille[69]) &&
(grille[64] != grille[70]) &&
(grille[64] != grille[71]) &&
(grille[65] != grille[66]) &&
(grille[65] != grille[67]) &&
(grille[65] != grille[68]) &&
(grille[65] != grille[69]) &&
(grille[65] != grille[70]) &&
(grille[65] != grille[71]) &&
(grille[66] != grille[67]) &&
(grille[66] != grille[68]) &&
(grille[66] != grille[69]) &&
(grille[66] != grille[70]) &&
(grille[66] != grille[71]) &&
(grille[67] != grille[68]) &&
(grille[67] != grille[69]) &&
(grille[67] != grille[70]) &&
(grille[67] != grille[71]) &&
(grille[68] != grille[69]) &&
(grille[68] != grille[70]) &&
(grille[68] != grille[71]) &&
(grille[69] != grille[70]) &&
(grille[69] != grille[71]) &&
(grille[70] != grille[71]) &&
(grille[72] != grille[73]) &&
(grille[72] != grille[74]) &&
(grille[72] != grille[75]) &&
(grille[72] != grille[76]) &&
(grille[72] != grille[77]) &&
(grille[72] != grille[78]) &&
(grille[72] != grille[79]) &&
(grille[72] != grille[80]) &&
(grille[73] != grille[74]) &&
(grille[73] != grille[75]) &&
(grille[73] != grille[76]) &&
(grille[73] != grille[77]) &&
(grille[73] != grille[78]) &&
(grille[73] != grille[79]) &&
(grille[73] != grille[80]) &&
(grille[74] != grille[75]) &&
(grille[74] != grille[76]) &&
(grille[74] != grille[77]) &&
(grille[74] != grille[78]) &&
(grille[74] != grille[79]) &&
(grille[74] != grille[80]) &&
(grille[75] != grille[76]) &&
(grille[75] != grille[77]) &&
(grille[75] != grille[78]) &&
(grille[75] != grille[79]) &&
(grille[75] != grille[80]) &&
(grille[76] != grille[77]) &&
(grille[76] != grille[78]) &&
(grille[76] != grille[79]) &&
(grille[76] != grille[80]) &&
(grille[77] != grille[78]) &&
(grille[77] != grille[79]) &&
(grille[77] != grille[80]) &&
(grille[78] != grille[79]) &&
(grille[78] != grille[80]) &&
(grille[79] != grille[80]) &&
(grille[0] != grille[9]) &&
(grille[0] != grille[18]) &&
(grille[0] != grille[27]) &&
(grille[0] != grille[36]) &&
(grille[0] != grille[45]) &&
(grille[0] != grille[54]) &&
(grille[0] != grille[63]) &&
(grille[0] != grille[72]) &&
(grille[9] != grille[18]) &&
(grille[9] != grille[27]) &&
(grille[9] != grille[36]) &&
(grille[9] != grille[45]) &&
(grille[9] != grille[54]) &&
(grille[9] != grille[63]) &&
(grille[9] != grille[72]) &&
(grille[18] != grille[27]) &&
(grille[18] != grille[36]) &&
(grille[18] != grille[45]) &&
(grille[18] != grille[54]) &&
(grille[18] != grille[63]) &&
(grille[18] != grille[72]) &&
(grille[27] != grille[36]) &&
(grille[27] != grille[45]) &&
(grille[27] != grille[54]) &&
(grille[27] != grille[63]) &&
(grille[27] != grille[72]) &&
(grille[36] != grille[45]) &&
(grille[36] != grille[54]) &&
(grille[36] != grille[63]) &&
(grille[36] != grille[72]) &&
(grille[45] != grille[54]) &&
(grille[45] != grille[63]) &&
(grille[45] != grille[72]) &&
(grille[54] != grille[63]) &&
(grille[54] != grille[72]) &&
(grille[63] != grille[72]) &&
(grille[1] != grille[10]) &&
(grille[1] != grille[19]) &&
(grille[1] != grille[28]) &&
(grille[1] != grille[37]) &&
(grille[1] != grille[46]) &&
(grille[1] != grille[55]) &&
(grille[1] != grille[64]) &&
(grille[1] != grille[73]) &&
(grille[10] != grille[19]) &&
(grille[10] != grille[28]) &&
(grille[10] != grille[37]) &&
(grille[10] != grille[46]) &&
(grille[10] != grille[55]) &&
(grille[10] != grille[64]) &&
(grille[10] != grille[73]) &&
(grille[19] != grille[28]) &&
(grille[19] != grille[37]) &&
(grille[19] != grille[46]) &&
(grille[19] != grille[55]) &&
(grille[19] != grille[64]) &&
(grille[19] != grille[73]) &&
(grille[28] != grille[37]) &&
(grille[28] != grille[46]) &&
(grille[28] != grille[55]) &&
(grille[28] != grille[64]) &&
(grille[28] != grille[73]) &&
(grille[37] != grille[46]) &&
(grille[37] != grille[55]) &&
(grille[37] != grille[64]) &&
(grille[37] != grille[73]) &&
(grille[46] != grille[55]) &&
(grille[46] != grille[64]) &&
(grille[46] != grille[73]) &&
(grille[55] != grille[64]) &&
(grille[55] != grille[73]) &&
(grille[64] != grille[73]) &&
(grille[2] != grille[11]) &&
(grille[2] != grille[20]) &&
(grille[2] != grille[29]) &&
(grille[2] != grille[38]) &&
(grille[2] != grille[47]) &&
(grille[2] != grille[56]) &&
(grille[2] != grille[65]) &&
(grille[2] != grille[74]) &&
(grille[11] != grille[20]) &&
(grille[11] != grille[29]) &&
(grille[11] != grille[38]) &&
(grille[11] != grille[47]) &&
(grille[11] != grille[56]) &&
(grille[11] != grille[65]) &&
(grille[11] != grille[74]) &&
(grille[20] != grille[29]) &&
(grille[20] != grille[38]) &&
(grille[20] != grille[47]) &&
(grille[20] != grille[56]) &&
(grille[20] != grille[65]) &&
(grille[20] != grille[74]) &&
(grille[29] != grille[38]) &&
(grille[29] != grille[47]) &&
(grille[29] != grille[56]) &&
(grille[29] != grille[65]) &&
(grille[29] != grille[74]) &&
(grille[38] != grille[47]) &&
(grille[38] != grille[56]) &&
(grille[38] != grille[65]) &&
(grille[38] != grille[74]) &&
(grille[47] != grille[56]) &&
(grille[47] != grille[65]) &&
(grille[47] != grille[74]) &&
(grille[56] != grille[65]) &&
(grille[56] != grille[74]) &&
(grille[65] != grille[74]) &&
(grille[3] != grille[12]) &&
(grille[3] != grille[21]) &&
(grille[3] != grille[30]) &&
(grille[3] != grille[39]) &&
(grille[3] != grille[48]) &&
(grille[3] != grille[57]) &&
(grille[3] != grille[66]) &&
(grille[3] != grille[75]) &&
(grille[12] != grille[21]) &&
(grille[12] != grille[30]) &&
(grille[12] != grille[39]) &&
(grille[12] != grille[48]) &&
(grille[12] != grille[57]) &&
(grille[12] != grille[66]) &&
(grille[12] != grille[75]) &&
(grille[21] != grille[30]) &&
(grille[21] != grille[39]) &&
(grille[21] != grille[48]) &&
(grille[21] != grille[57]) &&
(grille[21] != grille[66]) &&
(grille[21] != grille[75]) &&
(grille[30] != grille[39]) &&
(grille[30] != grille[48]) &&
(grille[30] != grille[57]) &&
(grille[30] != grille[66]) &&
(grille[30] != grille[75]) &&
(grille[39] != grille[48]) &&
(grille[39] != grille[57]) &&
(grille[39] != grille[66]) &&
(grille[39] != grille[75]) &&
(grille[48] != grille[57]) &&
(grille[48] != grille[66]) &&
(grille[48] != grille[75]) &&
(grille[57] != grille[66]) &&
(grille[57] != grille[75]) &&
(grille[66] != grille[75]) &&
(grille[4] != grille[13]) &&
(grille[4] != grille[22]) &&
(grille[4] != grille[31]) &&
(grille[4] != grille[40]) &&
(grille[4] != grille[49]) &&
(grille[4] != grille[58]) &&
(grille[4] != grille[67]) &&
(grille[4] != grille[76]) &&
(grille[13] != grille[22]) &&
(grille[13] != grille[31]) &&
(grille[13] != grille[40]) &&
(grille[13] != grille[49]) &&
(grille[13] != grille[58]) &&
(grille[13] != grille[67]) &&
(grille[13] != grille[76]) &&
(grille[22] != grille[31]) &&
(grille[22] != grille[40]) &&
(grille[22] != grille[49]) &&
(grille[22] != grille[58]) &&
(grille[22] != grille[67]) &&
(grille[22] != grille[76]) &&
(grille[31] != grille[40]) &&
(grille[31] != grille[49]) &&
(grille[31] != grille[58]) &&
(grille[31] != grille[67]) &&
(grille[31] != grille[76]) &&
(grille[40] != grille[49]) &&
(grille[40] != grille[58]) &&
(grille[40] != grille[67]) &&
(grille[40] != grille[76]) &&
(grille[49] != grille[58]) &&
(grille[49] != grille[67]) &&
(grille[49] != grille[76]) &&
(grille[58] != grille[67]) &&
(grille[58] != grille[76]) &&
(grille[67] != grille[76]) &&
(grille[5] != grille[14]) &&
(grille[5] != grille[23]) &&
(grille[5] != grille[32]) &&
(grille[5] != grille[41]) &&
(grille[5] != grille[50]) &&
(grille[5] != grille[59]) &&
(grille[5] != grille[68]) &&
(grille[5] != grille[77]) &&
(grille[14] != grille[23]) &&
(grille[14] != grille[32]) &&
(grille[14] != grille[41]) &&
(grille[14] != grille[50]) &&
(grille[14] != grille[59]) &&
(grille[14] != grille[68]) &&
(grille[14] != grille[77]) &&
(grille[23] != grille[32]) &&
(grille[23] != grille[41]) &&
(grille[23] != grille[50]) &&
(grille[23] != grille[59]) &&
(grille[23] != grille[68]) &&
(grille[23] != grille[77]) &&
(grille[32] != grille[41]) &&
(grille[32] != grille[50]) &&
(grille[32] != grille[59]) &&
(grille[32] != grille[68]) &&
(grille[32] != grille[77]) &&
(grille[41] != grille[50]) &&
(grille[41] != grille[59]) &&
(grille[41] != grille[68]) &&
(grille[41] != grille[77]) &&
(grille[50] != grille[59]) &&
(grille[50] != grille[68]) &&
(grille[50] != grille[77]) &&
(grille[59] != grille[68]) &&
(grille[59] != grille[77]) &&
(grille[68] != grille[77]) &&
(grille[6] != grille[15]) &&
(grille[6] != grille[24]) &&
(grille[6] != grille[33]) &&
(grille[6] != grille[42]) &&
(grille[6] != grille[51]) &&
(grille[6] != grille[60]) &&
(grille[6] != grille[69]) &&
(grille[6] != grille[78]) &&
(grille[15] != grille[24]) &&
(grille[15] != grille[33]) &&
(grille[15] != grille[42]) &&
(grille[15] != grille[51]) &&
(grille[15] != grille[60]) &&
(grille[15] != grille[69]) &&
(grille[15] != grille[78]) &&
(grille[24] != grille[33]) &&
(grille[24] != grille[42]) &&
(grille[24] != grille[51]) &&
(grille[24] != grille[60]) &&
(grille[24] != grille[69]) &&
(grille[24] != grille[78]) &&
(grille[33] != grille[42]) &&
(grille[33] != grille[51]) &&
(grille[33] != grille[60]) &&
(grille[33] != grille[69]) &&
(grille[33] != grille[78]) &&
(grille[42] != grille[51]) &&
(grille[42] != grille[60]) &&
(grille[42] != grille[69]) &&
(grille[42] != grille[78]) &&
(grille[51] != grille[60]) &&
(grille[51] != grille[69]) &&
(grille[51] != grille[78]) &&
(grille[60] != grille[69]) &&
(grille[60] != grille[78]) &&
(grille[69] != grille[78]) &&
(grille[7] != grille[16]) &&
(grille[7] != grille[25]) &&
(grille[7] != grille[34]) &&
(grille[7] != grille[43]) &&
(grille[7] != grille[52]) &&
(grille[7] != grille[61]) &&
(grille[7] != grille[70]) &&
(grille[7] != grille[79]) &&
(grille[16] != grille[25]) &&
(grille[16] != grille[34]) &&
(grille[16] != grille[43]) &&
(grille[16] != grille[52]) &&
(grille[16] != grille[61]) &&
(grille[16] != grille[70]) &&
(grille[16] != grille[79]) &&
(grille[25] != grille[34]) &&
(grille[25] != grille[43]) &&
(grille[25] != grille[52]) &&
(grille[25] != grille[61]) &&
(grille[25] != grille[70]) &&
(grille[25] != grille[79]) &&
(grille[34] != grille[43]) &&
(grille[34] != grille[52]) &&
(grille[34] != grille[61]) &&
(grille[34] != grille[70]) &&
(grille[34] != grille[79]) &&
(grille[43] != grille[52]) &&
(grille[43] != grille[61]) &&
(grille[43] != grille[70]) &&
(grille[43] != grille[79]) &&
(grille[52] != grille[61]) &&
(grille[52] != grille[70]) &&
(grille[52] != grille[79]) &&
(grille[61] != grille[70]) &&
(grille[61] != grille[79]) &&
(grille[70] != grille[79]) &&
(grille[8] != grille[17]) &&
(grille[8] != grille[26]) &&
(grille[8] != grille[35]) &&
(grille[8] != grille[44]) &&
(grille[8] != grille[53]) &&
(grille[8] != grille[62]) &&
(grille[8] != grille[71]) &&
(grille[8] != grille[80]) &&
(grille[17] != grille[26]) &&
(grille[17] != grille[35]) &&
(grille[17] != grille[44]) &&
(grille[17] != grille[53]) &&
(grille[17] != grille[62]) &&
(grille[17] != grille[71]) &&
(grille[17] != grille[80]) &&
(grille[26] != grille[35]) &&
(grille[26] != grille[44]) &&
(grille[26] != grille[53]) &&
(grille[26] != grille[62]) &&
(grille[26] != grille[71]) &&
(grille[26] != grille[80]) &&
(grille[35] != grille[44]) &&
(grille[35] != grille[53]) &&
(grille[35] != grille[62]) &&
(grille[35] != grille[71]) &&
(grille[35] != grille[80]) &&
(grille[44] != grille[53]) &&
(grille[44] != grille[62]) &&
(grille[44] != grille[71]) &&
(grille[44] != grille[80]) &&
(grille[53] != grille[62]) &&
(grille[53] != grille[71]) &&
(grille[53] != grille[80]) &&
(grille[62] != grille[71]) &&
(grille[62] != grille[80]) &&
(grille[71] != grille[80]) &&
(grille[0] != grille[1]) &&
(grille[0] != grille[2]) &&
(grille[0] != grille[9]) &&
(grille[0] != grille[10]) &&
(grille[0] != grille[11]) &&
(grille[0] != grille[18]) &&
(grille[0] != grille[19]) &&
(grille[0] != grille[20]) &&
(grille[1] != grille[0]) &&
(grille[1] != grille[2]) &&
(grille[1] != grille[9]) &&
(grille[1] != grille[10]) &&
(grille[1] != grille[11]) &&
(grille[1] != grille[18]) &&
(grille[1] != grille[19]) &&
(grille[1] != grille[20]) &&
(grille[2] != grille[0]) &&
(grille[2] != grille[1]) &&
(grille[2] != grille[9]) &&
(grille[2] != grille[10]) &&
(grille[2] != grille[11]) &&
(grille[2] != grille[18]) &&
(grille[2] != grille[19]) &&
(grille[2] != grille[20]) &&
(grille[9] != grille[0]) &&
(grille[9] != grille[1]) &&
(grille[9] != grille[2]) &&
(grille[9] != grille[10]) &&
(grille[9] != grille[11]) &&
(grille[9] != grille[18]) &&
(grille[9] != grille[19]) &&
(grille[9] != grille[20]) &&
(grille[10] != grille[0]) &&
(grille[10] != grille[1]) &&
(grille[10] != grille[2]) &&
(grille[10] != grille[9]) &&
(grille[10] != grille[11]) &&
(grille[10] != grille[18]) &&
(grille[10] != grille[19]) &&
(grille[10] != grille[20]) &&
(grille[11] != grille[0]) &&
(grille[11] != grille[1]) &&
(grille[11] != grille[2]) &&
(grille[11] != grille[9]) &&
(grille[11] != grille[10]) &&
(grille[11] != grille[18]) &&
(grille[11] != grille[19]) &&
(grille[11] != grille[20]) &&
(grille[18] != grille[0]) &&
(grille[18] != grille[1]) &&
(grille[18] != grille[2]) &&
(grille[18] != grille[9]) &&
(grille[18] != grille[10]) &&
(grille[18] != grille[11]) &&
(grille[18] != grille[19]) &&
(grille[18] != grille[20]) &&
(grille[19] != grille[0]) &&
(grille[19] != grille[1]) &&
(grille[19] != grille[2]) &&
(grille[19] != grille[9]) &&
(grille[19] != grille[10]) &&
(grille[19] != grille[11]) &&
(grille[19] != grille[18]) &&
(grille[19] != grille[20]) &&
(grille[20] != grille[0]) &&
(grille[20] != grille[1]) &&
(grille[20] != grille[2]) &&
(grille[20] != grille[9]) &&
(grille[20] != grille[10]) &&
(grille[20] != grille[11]) &&
(grille[20] != grille[18]) &&
(grille[20] != grille[19]) &&
(grille[3] != grille[4]) &&
(grille[3] != grille[5]) &&
(grille[3] != grille[12]) &&
(grille[3] != grille[13]) &&
(grille[3] != grille[14]) &&
(grille[3] != grille[21]) &&
(grille[3] != grille[22]) &&
(grille[3] != grille[23]) &&
(grille[4] != grille[3]) &&
(grille[4] != grille[5]) &&
(grille[4] != grille[12]) &&
(grille[4] != grille[13]) &&
(grille[4] != grille[14]) &&
(grille[4] != grille[21]) &&
(grille[4] != grille[22]) &&
(grille[4] != grille[23]) &&
(grille[5] != grille[3]) &&
(grille[5] != grille[4]) &&
(grille[5] != grille[12]) &&
(grille[5] != grille[13]) &&
(grille[5] != grille[14]) &&
(grille[5] != grille[21]) &&
(grille[5] != grille[22]) &&
(grille[5] != grille[23]) &&
(grille[12] != grille[3]) &&
(grille[12] != grille[4]) &&
(grille[12] != grille[5]) &&
(grille[12] != grille[13]) &&
(grille[12] != grille[14]) &&
(grille[12] != grille[21]) &&
(grille[12] != grille[22]) &&
(grille[12] != grille[23]) &&
(grille[13] != grille[3]) &&
(grille[13] != grille[4]) &&
(grille[13] != grille[5]) &&
(grille[13] != grille[12]) &&
(grille[13] != grille[14]) &&
(grille[13] != grille[21]) &&
(grille[13] != grille[22]) &&
(grille[13] != grille[23]) &&
(grille[14] != grille[3]) &&
(grille[14] != grille[4]) &&
(grille[14] != grille[5]) &&
(grille[14] != grille[12]) &&
(grille[14] != grille[13]) &&
(grille[14] != grille[21]) &&
(grille[14] != grille[22]) &&
(grille[14] != grille[23]) &&
(grille[21] != grille[3]) &&
(grille[21] != grille[4]) &&
(grille[21] != grille[5]) &&
(grille[21] != grille[12]) &&
(grille[21] != grille[13]) &&
(grille[21] != grille[14]) &&
(grille[21] != grille[22]) &&
(grille[21] != grille[23]) &&
(grille[22] != grille[3]) &&
(grille[22] != grille[4]) &&
(grille[22] != grille[5]) &&
(grille[22] != grille[12]) &&
(grille[22] != grille[13]) &&
(grille[22] != grille[14]) &&
(grille[22] != grille[21]) &&
(grille[22] != grille[23]) &&
(grille[23] != grille[3]) &&
(grille[23] != grille[4]) &&
(grille[23] != grille[5]) &&
(grille[23] != grille[12]) &&
(grille[23] != grille[13]) &&
(grille[23] != grille[14]) &&
(grille[23] != grille[21]) &&
(grille[23] != grille[22]) &&
(grille[6] != grille[7]) &&
(grille[6] != grille[8]) &&
(grille[6] != grille[15]) &&
(grille[6] != grille[16]) &&
(grille[6] != grille[17]) &&
(grille[6] != grille[24]) &&
(grille[6] != grille[25]) &&
(grille[6] != grille[26]) &&
(grille[7] != grille[6]) &&
(grille[7] != grille[8]) &&
(grille[7] != grille[15]) &&
(grille[7] != grille[16]) &&
(grille[7] != grille[17]) &&
(grille[7] != grille[24]) &&
(grille[7] != grille[25]) &&
(grille[7] != grille[26]) &&
(grille[8] != grille[6]) &&
(grille[8] != grille[7]) &&
(grille[8] != grille[15]) &&
(grille[8] != grille[16]) &&
(grille[8] != grille[17]) &&
(grille[8] != grille[24]) &&
(grille[8] != grille[25]) &&
(grille[8] != grille[26]) &&
(grille[15] != grille[6]) &&
(grille[15] != grille[7]) &&
(grille[15] != grille[8]) &&
(grille[15] != grille[16]) &&
(grille[15] != grille[17]) &&
(grille[15] != grille[24]) &&
(grille[15] != grille[25]) &&
(grille[15] != grille[26]) &&
(grille[16] != grille[6]) &&
(grille[16] != grille[7]) &&
(grille[16] != grille[8]) &&
(grille[16] != grille[15]) &&
(grille[16] != grille[17]) &&
(grille[16] != grille[24]) &&
(grille[16] != grille[25]) &&
(grille[16] != grille[26]) &&
(grille[17] != grille[6]) &&
(grille[17] != grille[7]) &&
(grille[17] != grille[8]) &&
(grille[17] != grille[15]) &&
(grille[17] != grille[16]) &&
(grille[17] != grille[24]) &&
(grille[17] != grille[25]) &&
(grille[17] != grille[26]) &&
(grille[24] != grille[6]) &&
(grille[24] != grille[7]) &&
(grille[24] != grille[8]) &&
(grille[24] != grille[15]) &&
(grille[24] != grille[16]) &&
(grille[24] != grille[17]) &&
(grille[24] != grille[25]) &&
(grille[24] != grille[26]) &&
(grille[25] != grille[6]) &&
(grille[25] != grille[7]) &&
(grille[25] != grille[8]) &&
(grille[25] != grille[15]) &&
(grille[25] != grille[16]) &&
(grille[25] != grille[17]) &&
(grille[25] != grille[24]) &&
(grille[25] != grille[26]) &&
(grille[26] != grille[6]) &&
(grille[26] != grille[7]) &&
(grille[26] != grille[8]) &&
(grille[26] != grille[15]) &&
(grille[26] != grille[16]) &&
(grille[26] != grille[17]) &&
(grille[26] != grille[24]) &&
(grille[26] != grille[25]) &&
(grille[27] != grille[28]) &&
(grille[27] != grille[29]) &&
(grille[27] != grille[36]) &&
(grille[27] != grille[37]) &&
(grille[27] != grille[38]) &&
(grille[27] != grille[45]) &&
(grille[27] != grille[46]) &&
(grille[27] != grille[47]) &&
(grille[28] != grille[27]) &&
(grille[28] != grille[29]) &&
(grille[28] != grille[36]) &&
(grille[28] != grille[37]) &&
(grille[28] != grille[38]) &&
(grille[28] != grille[45]) &&
(grille[28] != grille[46]) &&
(grille[28] != grille[47]) &&
(grille[29] != grille[27]) &&
(grille[29] != grille[28]) &&
(grille[29] != grille[36]) &&
(grille[29] != grille[37]) &&
(grille[29] != grille[38]) &&
(grille[29] != grille[45]) &&
(grille[29] != grille[46]) &&
(grille[29] != grille[47]) &&
(grille[36] != grille[27]) &&
(grille[36] != grille[28]) &&
(grille[36] != grille[29]) &&
(grille[36] != grille[37]) &&
(grille[36] != grille[38]) &&
(grille[36] != grille[45]) &&
(grille[36] != grille[46]) &&
(grille[36] != grille[47]) &&
(grille[37] != grille[27]) &&
(grille[37] != grille[28]) &&
(grille[37] != grille[29]) &&
(grille[37] != grille[36]) &&
(grille[37] != grille[38]) &&
(grille[37] != grille[45]) &&
(grille[37] != grille[46]) &&
(grille[37] != grille[47]) &&
(grille[38] != grille[27]) &&
(grille[38] != grille[28]) &&
(grille[38] != grille[29]) &&
(grille[38] != grille[36]) &&
(grille[38] != grille[37]) &&
(grille[38] != grille[45]) &&
(grille[38] != grille[46]) &&
(grille[38] != grille[47]) &&
(grille[45] != grille[27]) &&
(grille[45] != grille[28]) &&
(grille[45] != grille[29]) &&
(grille[45] != grille[36]) &&
(grille[45] != grille[37]) &&
(grille[45] != grille[38]) &&
(grille[45] != grille[46]) &&
(grille[45] != grille[47]) &&
(grille[46] != grille[27]) &&
(grille[46] != grille[28]) &&
(grille[46] != grille[29]) &&
(grille[46] != grille[36]) &&
(grille[46] != grille[37]) &&
(grille[46] != grille[38]) &&
(grille[46] != grille[45]) &&
(grille[46] != grille[47]) &&
(grille[47] != grille[27]) &&
(grille[47] != grille[28]) &&
(grille[47] != grille[29]) &&
(grille[47] != grille[36]) &&
(grille[47] != grille[37]) &&
(grille[47] != grille[38]) &&
(grille[47] != grille[45]) &&
(grille[47] != grille[46]) &&
(grille[30] != grille[31]) &&
(grille[30] != grille[32]) &&
(grille[30] != grille[39]) &&
(grille[30] != grille[40]) &&
(grille[30] != grille[41]) &&
(grille[30] != grille[48]) &&
(grille[30] != grille[49]) &&
(grille[30] != grille[50]) &&
(grille[31] != grille[30]) &&
(grille[31] != grille[32]) &&
(grille[31] != grille[39]) &&
(grille[31] != grille[40]) &&
(grille[31] != grille[41]) &&
(grille[31] != grille[48]) &&
(grille[31] != grille[49]) &&
(grille[31] != grille[50]) &&
(grille[32] != grille[30]) &&
(grille[32] != grille[31]) &&
(grille[32] != grille[39]) &&
(grille[32] != grille[40]) &&
(grille[32] != grille[41]) &&
(grille[32] != grille[48]) &&
(grille[32] != grille[49]) &&
(grille[32] != grille[50]) &&
(grille[39] != grille[30]) &&
(grille[39] != grille[31]) &&
(grille[39] != grille[32]) &&
(grille[39] != grille[40]) &&
(grille[39] != grille[41]) &&
(grille[39] != grille[48]) &&
(grille[39] != grille[49]) &&
(grille[39] != grille[50]) &&
(grille[40] != grille[30]) &&
(grille[40] != grille[31]) &&
(grille[40] != grille[32]) &&
(grille[40] != grille[39]) &&
(grille[40] != grille[41]) &&
(grille[40] != grille[48]) &&
(grille[40] != grille[49]) &&
(grille[40] != grille[50]) &&
(grille[41] != grille[30]) &&
(grille[41] != grille[31]) &&
(grille[41] != grille[32]) &&
(grille[41] != grille[39]) &&
(grille[41] != grille[40]) &&
(grille[41] != grille[48]) &&
(grille[41] != grille[49]) &&
(grille[41] != grille[50]) &&
(grille[48] != grille[30]) &&
(grille[48] != grille[31]) &&
(grille[48] != grille[32]) &&
(grille[48] != grille[39]) &&
(grille[48] != grille[40]) &&
(grille[48] != grille[41]) &&
(grille[48] != grille[49]) &&
(grille[48] != grille[50]) &&
(grille[49] != grille[30]) &&
(grille[49] != grille[31]) &&
(grille[49] != grille[32]) &&
(grille[49] != grille[39]) &&
(grille[49] != grille[40]) &&
(grille[49] != grille[41]) &&
(grille[49] != grille[48]) &&
(grille[49] != grille[50]) &&
(grille[50] != grille[30]) &&
(grille[50] != grille[31]) &&
(grille[50] != grille[32]) &&
(grille[50] != grille[39]) &&
(grille[50] != grille[40]) &&
(grille[50] != grille[41]) &&
(grille[50] != grille[48]) &&
(grille[50] != grille[49]) &&
(grille[33] != grille[34]) &&
(grille[33] != grille[35]) &&
(grille[33] != grille[42]) &&
(grille[33] != grille[43]) &&
(grille[33] != grille[44]) &&
(grille[33] != grille[51]) &&
(grille[33] != grille[52]) &&
(grille[33] != grille[53]) &&
(grille[34] != grille[33]) &&
(grille[34] != grille[35]) &&
(grille[34] != grille[42]) &&
(grille[34] != grille[43]) &&
(grille[34] != grille[44]) &&
(grille[34] != grille[51]) &&
(grille[34] != grille[52]) &&
(grille[34] != grille[53]) &&
(grille[35] != grille[33]) &&
(grille[35] != grille[34]) &&
(grille[35] != grille[42]) &&
(grille[35] != grille[43]) &&
(grille[35] != grille[44]) &&
(grille[35] != grille[51]) &&
(grille[35] != grille[52]) &&
(grille[35] != grille[53]) &&
(grille[42] != grille[33]) &&
(grille[42] != grille[34]) &&
(grille[42] != grille[35]) &&
(grille[42] != grille[43]) &&
(grille[42] != grille[44]) &&
(grille[42] != grille[51]) &&
(grille[42] != grille[52]) &&
(grille[42] != grille[53]) &&
(grille[43] != grille[33]) &&
(grille[43] != grille[34]) &&
(grille[43] != grille[35]) &&
(grille[43] != grille[42]) &&
(grille[43] != grille[44]) &&
(grille[43] != grille[51]) &&
(grille[43] != grille[52]) &&
(grille[43] != grille[53]) &&
(grille[44] != grille[33]) &&
(grille[44] != grille[34]) &&
(grille[44] != grille[35]) &&
(grille[44] != grille[42]) &&
(grille[44] != grille[43]) &&
(grille[44] != grille[51]) &&
(grille[44] != grille[52]) &&
(grille[44] != grille[53]) &&
(grille[51] != grille[33]) &&
(grille[51] != grille[34]) &&
(grille[51] != grille[35]) &&
(grille[51] != grille[42]) &&
(grille[51] != grille[43]) &&
(grille[51] != grille[44]) &&
(grille[51] != grille[52]) &&
(grille[51] != grille[53]) &&
(grille[52] != grille[33]) &&
(grille[52] != grille[34]) &&
(grille[52] != grille[35]) &&
(grille[52] != grille[42]) &&
(grille[52] != grille[43]) &&
(grille[52] != grille[44]) &&
(grille[52] != grille[51]) &&
(grille[52] != grille[53]) &&
(grille[53] != grille[33]) &&
(grille[53] != grille[34]) &&
(grille[53] != grille[35]) &&
(grille[53] != grille[42]) &&
(grille[53] != grille[43]) &&
(grille[53] != grille[44]) &&
(grille[53] != grille[51]) &&
(grille[53] != grille[52]) &&
(grille[54] != grille[55]) &&
(grille[54] != grille[56]) &&
(grille[54] != grille[63]) &&
(grille[54] != grille[64]) &&
(grille[54] != grille[65]) &&
(grille[54] != grille[72]) &&
(grille[54] != grille[73]) &&
(grille[54] != grille[74]) &&
(grille[55] != grille[54]) &&
(grille[55] != grille[56]) &&
(grille[55] != grille[63]) &&
(grille[55] != grille[64]) &&
(grille[55] != grille[65]) &&
(grille[55] != grille[72]) &&
(grille[55] != grille[73]) &&
(grille[55] != grille[74]) &&
(grille[56] != grille[54]) &&
(grille[56] != grille[55]) &&
(grille[56] != grille[63]) &&
(grille[56] != grille[64]) &&
(grille[56] != grille[65]) &&
(grille[56] != grille[72]) &&
(grille[56] != grille[73]) &&
(grille[56] != grille[74]) &&
(grille[63] != grille[54]) &&
(grille[63] != grille[55]) &&
(grille[63] != grille[56]) &&
(grille[63] != grille[64]) &&
(grille[63] != grille[65]) &&
(grille[63] != grille[72]) &&
(grille[63] != grille[73]) &&
(grille[63] != grille[74]) &&
(grille[64] != grille[54]) &&
(grille[64] != grille[55]) &&
(grille[64] != grille[56]) &&
(grille[64] != grille[63]) &&
(grille[64] != grille[65]) &&
(grille[64] != grille[72]) &&
(grille[64] != grille[73]) &&
(grille[64] != grille[74]) &&
(grille[65] != grille[54]) &&
(grille[65] != grille[55]) &&
(grille[65] != grille[56]) &&
(grille[65] != grille[63]) &&
(grille[65] != grille[64]) &&
(grille[65] != grille[72]) &&
(grille[65] != grille[73]) &&
(grille[65] != grille[74]) &&
(grille[72] != grille[54]) &&
(grille[72] != grille[55]) &&
(grille[72] != grille[56]) &&
(grille[72] != grille[63]) &&
(grille[72] != grille[64]) &&
(grille[72] != grille[65]) &&
(grille[72] != grille[73]) &&
(grille[72] != grille[74]) &&
(grille[73] != grille[54]) &&
(grille[73] != grille[55]) &&
(grille[73] != grille[56]) &&
(grille[73] != grille[63]) &&
(grille[73] != grille[64]) &&
(grille[73] != grille[65]) &&
(grille[73] != grille[72]) &&
(grille[73] != grille[74]) &&
(grille[74] != grille[54]) &&
(grille[74] != grille[55]) &&
(grille[74] != grille[56]) &&
(grille[74] != grille[63]) &&
(grille[74] != grille[64]) &&
(grille[74] != grille[65]) &&
(grille[74] != grille[72]) &&
(grille[74] != grille[73]) &&
(grille[57] != grille[58]) &&
(grille[57] != grille[59]) &&
(grille[57] != grille[66]) &&
(grille[57] != grille[67]) &&
(grille[57] != grille[68]) &&
(grille[57] != grille[75]) &&
(grille[57] != grille[76]) &&
(grille[57] != grille[77]) &&
(grille[58] != grille[57]) &&
(grille[58] != grille[59]) &&
(grille[58] != grille[66]) &&
(grille[58] != grille[67]) &&
(grille[58] != grille[68]) &&
(grille[58] != grille[75]) &&
(grille[58] != grille[76]) &&
(grille[58] != grille[77]) &&
(grille[59] != grille[57]) &&
(grille[59] != grille[58]) &&
(grille[59] != grille[66]) &&
(grille[59] != grille[67]) &&
(grille[59] != grille[68]) &&
(grille[59] != grille[75]) &&
(grille[59] != grille[76]) &&
(grille[59] != grille[77]) &&
(grille[66] != grille[57]) &&
(grille[66] != grille[58]) &&
(grille[66] != grille[59]) &&
(grille[66] != grille[67]) &&
(grille[66] != grille[68]) &&
(grille[66] != grille[75]) &&
(grille[66] != grille[76]) &&
(grille[66] != grille[77]) &&
(grille[67] != grille[57]) &&
(grille[67] != grille[58]) &&
(grille[67] != grille[59]) &&
(grille[67] != grille[66]) &&
(grille[67] != grille[68]) &&
(grille[67] != grille[75]) &&
(grille[67] != grille[76]) &&
(grille[67] != grille[77]) &&
(grille[68] != grille[57]) &&
(grille[68] != grille[58]) &&
(grille[68] != grille[59]) &&
(grille[68] != grille[66]) &&
(grille[68] != grille[67]) &&
(grille[68] != grille[75]) &&
(grille[68] != grille[76]) &&
(grille[68] != grille[77]) &&
(grille[75] != grille[57]) &&
(grille[75] != grille[58]) &&
(grille[75] != grille[59]) &&
(grille[75] != grille[66]) &&
(grille[75] != grille[67]) &&
(grille[75] != grille[68]) &&
(grille[75] != grille[76]) &&
(grille[75] != grille[77]) &&
(grille[76] != grille[57]) &&
(grille[76] != grille[58]) &&
(grille[76] != grille[59]) &&
(grille[76] != grille[66]) &&
(grille[76] != grille[67]) &&
(grille[76] != grille[68]) &&
(grille[76] != grille[75]) &&
(grille[76] != grille[77]) &&
(grille[77] != grille[57]) &&
(grille[77] != grille[58]) &&
(grille[77] != grille[59]) &&
(grille[77] != grille[66]) &&
(grille[77] != grille[67]) &&
(grille[77] != grille[68]) &&
(grille[77] != grille[75]) &&
(grille[77] != grille[76]) &&
(grille[60] != grille[61]) &&
(grille[60] != grille[62]) &&
(grille[60] != grille[69]) &&
(grille[60] != grille[70]) &&
(grille[60] != grille[71]) &&
(grille[60] != grille[78]) &&
(grille[60] != grille[79]) &&
(grille[60] != grille[80]) &&
(grille[61] != grille[60]) &&
(grille[61] != grille[62]) &&
(grille[61] != grille[69]) &&
(grille[61] != grille[70]) &&
(grille[61] != grille[71]) &&
(grille[61] != grille[78]) &&
(grille[61] != grille[79]) &&
(grille[61] != grille[80]) &&
(grille[62] != grille[60]) &&
(grille[62] != grille[61]) &&
(grille[62] != grille[69]) &&
(grille[62] != grille[70]) &&
(grille[62] != grille[71]) &&
(grille[62] != grille[78]) &&
(grille[62] != grille[79]) &&
(grille[62] != grille[80]) &&
(grille[69] != grille[60]) &&
(grille[69] != grille[61]) &&
(grille[69] != grille[62]) &&
(grille[69] != grille[70]) &&
(grille[69] != grille[71]) &&
(grille[69] != grille[78]) &&
(grille[69] != grille[79]) &&
(grille[69] != grille[80]) &&
(grille[70] != grille[60]) &&
(grille[70] != grille[61]) &&
(grille[70] != grille[62]) &&
(grille[70] != grille[69]) &&
(grille[70] != grille[71]) &&
(grille[70] != grille[78]) &&
(grille[70] != grille[79]) &&
(grille[70] != grille[80]) &&
(grille[71] != grille[60]) &&
(grille[71] != grille[61]) &&
(grille[71] != grille[62]) &&
(grille[71] != grille[69]) &&
(grille[71] != grille[70]) &&
(grille[71] != grille[78]) &&
(grille[71] != grille[79]) &&
(grille[71] != grille[80]) &&
(grille[78] != grille[60]) &&
(grille[78] != grille[61]) &&
(grille[78] != grille[62]) &&
(grille[78] != grille[69]) &&
(grille[78] != grille[70]) &&
(grille[78] != grille[71]) &&
(grille[78] != grille[79]) &&
(grille[78] != grille[80]) &&
(grille[79] != grille[60]) &&
(grille[79] != grille[61]) &&
(grille[79] != grille[62]) &&
(grille[79] != grille[69]) &&
(grille[79] != grille[70]) &&
(grille[79] != grille[71]) &&
(grille[79] != grille[78]) &&
(grille[79] != grille[80]) &&
(grille[80] != grille[60]) &&
(grille[80] != grille[61]) &&
(grille[80] != grille[62]) &&
(grille[80] != grille[69]) &&
(grille[80] != grille[70]) &&
(grille[80] != grille[71]) &&
(grille[80] != grille[78]) &&
(grille[80] != grille[79]) &&
(forall g:int in 0..80 { (0 < grille[g]) && (grille[g] <= 9) });
}
}